** Profile: "SCHEMATIC1-slewnew"  [ C:\ORCAD\ORCAD_16.6_LITE\TOOLS\CAPTURE\johnie -PSpiceFiles\SCHEMATIC1\slewnew.sim ] 

** Creating circuit file "slewnew.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/ORCAD/ORCAD_16.6_LITE/TOOLS/pspice/library/mosfets.lib" 
* From [PSPICE NETLIST] section of C:\Users\DELLGR\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10us 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
